*2 input Xor 1 output
 .include sky130nm.lib
 .option scale=10n
 Xxor2 neg_supply bin01 ain01 pos_supply xout_2_xor2 neg_supply pos_supply xor2
 Xxor2swap neg_supply ain01 bin01 pos_supply xout_2_swap_xor2 neg_supply pos_supply xor2
 Xxor3 neg_supply bin11 ain11 pos_supply xout_3_xor2 neg_supply pos_supply xor2
 Xxor3swap neg_supply ain11 bin11 pos_supply xout_3_swap_xor2 neg_supply pos_supply xor2

 *Xxor3 ain bin neg_supply neg_supply pos_supply pos_supply xoutmodel sky130_fd_sc_hd__xor2_1
 v3 pos_supply 0 1.0
 *v3 pos_supply 0 SINE(0 1.8 10000000 0 0 0)
 v4 neg_supply 0 0.0
 v2 ain01 0 PULSE 0.0 1.8 1n 20p 20p 2n 4ns
 v5 bin01 0 PULSE 0 1.8 1n 20p 20p 2n 4ns
 v6 ain11 0 PULSE 1.8 0.0 1n 20p 20p 2n 4ns
 v7 bin11 0 PULSE 1.8 0.0 1n 20p 20p 2n 4ns
.control  
 tran 1ps 50ns
 *plot  
 gnuplot gp v(ain01) v(bin01) v(xout_2_xor2)+2 v(xout_2_swap_xor2)+4 v(pos_supply)
 gnuplot gpa v(ain11) v(bin11) v(xout_3_xor2)+2 v(xout_3_swap_xor2)+4 v(pos_supply)
.endc
 
 
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 a_35_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=65 l=15
X1 VGND B a_35_297# VNB sky130_fd_pr__nfet_01v8 w=65 l=15
X2 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 w=65 l=15
X3 a_285_297# B VPWR VPB sky130_fd_pr__pfet_01v8 w=100 l=15
X4 VPWR A a_285_297# VPB sky130_fd_pr__pfet_01v8 w=100 l=15
X5 a_35_297# B a_117_297# VPB sky130_fd_pr__pfet_01v8 w=100 l=15
X6 a_117_297# A VPWR VPB sky130_fd_pr__pfet_01v8 w=100 l=15
X7 a_285_47# B X VNB sky130_fd_pr__nfet_01v8 w=65 l=15
X8 a_285_297# a_35_297# X VPB sky130_fd_pr__pfet_01v8 w=100 l=15
X9 VGND A a_285_47# VNB sky130_fd_pr__nfet_01v8 w=65 l=15
.ends

 .subckt xor2 VNB B A VPWR X VGND VPB
X0 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X1 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X2 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X3 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X4 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X5 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X6 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X7 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X8 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X9 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X10 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X11 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X12 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X13 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X14 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X15 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X16 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
X17 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=100 l=15
X19 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=65 l=15
C0 VGND VNB 1.01fF
C1 VPB VNB 1.22fF
.ends

.subckt riedelxor2_cyclic ainput binside ycyclic powin gndin SUB
Xxor2_0 SUB ycyclic ainput powin binside gndin powin xor2
Xxor2_1 SUB ainput binside powin ycyclic gndin powin xor2
C0 powin SUB 1.22fF 
C1 gndin SUB 2.64fF
C2 powin SUB 2.50fF
C3 ycyclic SUB 1.54fF
C4 ainput SUB 2.71fF
C5 powin SUB 1.22fF
.ends

 